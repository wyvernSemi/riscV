// Block name: core
// And now for some register addresses...
`define CSR_LOCAL_ADDR                      32'h00000000
`define CSR_LOCAL_ADDR_INT                  0

`define CSR_SCRATCH_ADDR                     5'h00
`define CSR_SCRATCH_ADDR_INT                 0

