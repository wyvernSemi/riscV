// Block name: zicsr
// And now for some register addresses...
`define RV32_MSTATUS_ADDR                    12'h300
`define RV32_MSTATUS_ADDR_INT                768
`define RV32_MSTATUS_UIE                     0:0
`define RV32_MSTATUS_SIE                     1:1
`define RV32_MSTATUS_MIE                     3:3
`define RV32_MSTATUS_UPIE                    4:4
`define RV32_MSTATUS_SPIE                    5:5
`define RV32_MSTATUS_MPIE                    7:7
`define RV32_MSTATUS_SPP                     8:8
`define RV32_MSTATUS_MPP                     12:11
`define RV32_MSTATUS_FS                      14:13
`define RV32_MSTATUS_XS                      16:15
`define RV32_MSTATUS_MPRV                    17:17
`define RV32_MSTATUS_SUM                     18:18
`define RV32_MSTATUS_MXR                     19:19
`define RV32_MSTATUS_TVM                     20:20
`define RV32_MSTATUS_TW                      21:21
`define RV32_MSTATUS_TSR                     22:22
`define RV32_MSTATUS_SD                      31:31
`define RV32_MISA_ADDR                       12'h301
`define RV32_MISA_ADDR_INT                   769
`define RV32_MISA_EXTENSIONS                 25:0
`define RV32_MISA_MXL                        31:30
`define RV32_MIE_ADDR                        12'h304
`define RV32_MIE_ADDR_INT                    772
`define RV32_MIE_USIE                        0:0
`define RV32_MIE_SSIE                        1:1
`define RV32_MIE_MSIE                        3:3
`define RV32_MIE_UTIE                        4:4
`define RV32_MIE_STIE                        5:5
`define RV32_MIE_MTIE                        7:7
`define RV32_MIE_UEIE                        8:8
`define RV32_MIE_SEIE                        9:9
`define RV32_MIE_MEIE                        11:11
`define RV32_MTVEC_ADDR                      12'h305
`define RV32_MTVEC_ADDR_INT                  773
`define RV32_MTVEC_MODE                      1:0
`define RV32_MTVEC_BASE                      31:2
`define RV32_MCOUNTEREN_ADDR                 12'h306
`define RV32_MCOUNTEREN_ADDR_INT             774
`define RV32_MCOUNTINHIBIT_ADDR              12'h320
`define RV32_MCOUNTINHIBIT_ADDR_INT          800
`define RV32_MCOUNTINHIBIT_CY                0:0
`define RV32_MCOUNTINHIBIT_IR                2:2
`define RV32_MSCRATCH_ADDR                   12'h340
`define RV32_MSCRATCH_ADDR_INT               832
`define RV32_MEPC_ADDR                       12'h341
`define RV32_MEPC_ADDR_INT                   833
`define RV32_MCAUSE_ADDR                     12'h342
`define RV32_MCAUSE_ADDR_INT                 834
`define RV32_MCAUSE_CODE                     3:0
`define RV32_MCAUSE_INTERRUPT                31:31
`define RV32_MTVAL_ADDR                      12'h343
`define RV32_MTVAL_ADDR_INT                  835
`define RV32_MIP_ADDR                        12'h344
`define RV32_MIP_ADDR_INT                    836
`define RV32_MIP_USIP                        0:0
`define RV32_MIP_SSIP                        1:1
`define RV32_MIP_MSIP                        3:3
`define RV32_MIP_UTIP                        4:4
`define RV32_MIP_STIP                        5:5
`define RV32_MIP_MTIP                        7:7
`define RV32_MIP_UEIP                        8:8
`define RV32_MIP_SEIP                        9:9
`define RV32_MIP_MEIP                        11:11
`define RV32_MCYCLE_ADDR                     12'hB00
`define RV32_MCYCLE_ADDR_INT                 2816
`define RV32_MINSTRET_ADDR                   12'hB02
`define RV32_MINSTRET_ADDR_INT               2818
`define RV32_MCYCLEH_ADDR                    12'hB80
`define RV32_MCYCLEH_ADDR_INT                2944
`define RV32_MINSTRETH_ADDR                  12'hB82
`define RV32_MINSTRETH_ADDR_INT              2946
`define RV32_UCYCLE_ADDR                     12'hC00
`define RV32_UCYCLE_ADDR_INT                 3072
`define RV32_UTIME_ADDR                      12'hC01
`define RV32_UTIME_ADDR_INT                  3073
`define RV32_UINSTRET_ADDR                   12'hC02
`define RV32_UINSTRET_ADDR_INT               3074
`define RV32_UCYCLEH_ADDR                    12'hC80
`define RV32_UCYCLEH_ADDR_INT                3200
`define RV32_UTIMEH_ADDR                     12'hC81
`define RV32_UTIMEH_ADDR_INT                 3201
`define RV32_UINSTRETH_ADDR                  12'hC82
`define RV32_UINSTRETH_ADDR_INT              3202
`define RV32_MVENDOR_ADDR                    12'hF11
`define RV32_MVENDOR_ADDR_INT                3857
`define RV32_MARCHID_ADDR                    12'hF12
`define RV32_MARCHID_ADDR_INT                3858
`define RV32_MIMPID_ADDR                     12'hF13
`define RV32_MIMPID_ADDR_INT                 3859
`define RV32_MHARTID_ADDR                    12'hF14
`define RV32_MHARTID_ADDR_INT                3860
`define RV32_CLK_FREQ_MHZ_ADDR               12'hFFF
`define RV32_CLK_FREQ_MHZ_ADDR_INT           4095

