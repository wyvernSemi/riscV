// -----------------------------------------------------------------------------
//  Title      : RISC-V RV32I decoder
//  Project    : rv32_cpu
// -----------------------------------------------------------------------------
//  File       : rv32.vh
//  Author     : Simon Southwell
//  Created    : 2021-12-03
//  Standard   : Verilog 2001
// -----------------------------------------------------------------------------
//  Description:
//  This file defines the top level common definitions
// -----------------------------------------------------------------------------
//  Copyright (c) 2021 Simon Southwell
// -----------------------------------------------------------------------------
//
//  This is free software: you can redistribute it and/or modify
//  it under the terms of the GNU General Public License as published by
//  the Free Software Foundation, either version 3 of the License, or
//  (at your option) any later version.
//
//  It is distributed in the hope that it will be useful,
//  but WITHOUT ANY WARRANTY; without even the implied warranty of
//  MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE. See the
//  GNU General Public License for more details.
//
//  You should have received a copy of the GNU General Public License
//  along with this code. If not, see <http://www.gnu.org/licenses/>.
//
// -----------------------------------------------------------------------------

// Definition to select synchronous or asynchronous reset

`ifndef RESET
//`define RESET 
`define RESET or negedge reset_n
`endif